module power_globals;
supply1 VPWR;
supply0 VGND;
supply1 VPB;
supply0 VNB;
endmodule
